Read Rope Circuit Simulation With Resistive Flexible Sensors
.include ./params.inc
r1 1 2 20k 
rOutEQ 2 0 18667
vcc 1 0 DC 5 
.control
unset askquit
op
print V(2)
echo output test > outresult.data  $ start new file
wrdata outresult V(2)
quit
.endc
.end