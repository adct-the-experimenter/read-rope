Read Rope Circuit Simulation With Resistive Flexible Sensors
.include ./params.inc
r1 1 2 20k 
r2_limit 2 0 10k 
r2_flex 2 0 valBend1 
vcc 1 0 DC 5 
.control
unset askquit
op
print V(2)
echo output test > outresult.data  $ start new file
wrdata outresult V(2)
quit
.endc
.end